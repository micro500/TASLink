library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity main is
    Port ( CLK : in std_logic;
           RX : in std_logic;
           TX : out std_logic;
           btn : in  STD_LOGIC_VECTOR (3 downto 0);
           p1_latch : in  STD_LOGIC;
           p1_clock : in  STD_LOGIC;
           p1_d0 : out STD_LOGIC;
           p1_d1 : out STD_LOGIC;
           p2_latch : in std_logic;
           p2_clock : in std_logic;
           p2_d0 : out std_logic;
           p2_d1 : out std_logic;
           p1_d0_oe : out std_logic;
           p2_d0_oe : out std_logic;
           p1_d1_oe : out std_logic;
           p2_d1_oe : out std_logic;
           debug : out STD_LOGIC_VECTOR (3 downto 0);
           l: out STD_LOGIC_VECTOR(3 downto 0));
end main;

architecture Behavioral of main is
  component shift_register is
    Port ( latch : in  STD_LOGIC;
           clock : in  STD_LOGIC;
           din : in  STD_LOGIC_VECTOR (7 downto 0);
           dout : out  STD_LOGIC;
           sin : in STD_LOGIC;
           clk : in std_logic);
  end component;
  
  component filter is
    Port ( signal_in : in  STD_LOGIC;
           clk : in  STD_LOGIC;
           signal_out : out  STD_LOGIC);
  end component;
  
  component toggle is
    Port ( signal_in : in  STD_LOGIC;
           signal_out : out  STD_LOGIC);
  end component;
  
  component UART is
    Port ( rx_data_out : out STD_LOGIC_VECTOR (7 downto 0);
           rx_data_was_recieved : in STD_LOGIC;
           rx_byte_waiting : out STD_LOGIC;
           clk : in  STD_LOGIC;

           rx_in : in STD_LOGIC;
           tx_data_in : in STD_LOGIC_VECTOR (7 downto 0);
           tx_buffer_full : out STD_LOGIC;
           tx_write : in STD_LOGIC;
           tx_out : out STD_LOGIC);
  end component;
  
  component controller is
    Port ( console_clock : in  STD_LOGIC;
           console_latch : in  STD_LOGIC;
           console_io : in  STD_LOGIC;
           console_d0 : out  STD_LOGIC;
           console_d1 : out  STD_LOGIC;
           console_d0_oe : out  STD_LOGIC;
           console_d1_oe : out  STD_LOGIC;
           data : in  STD_LOGIC_VECTOR (31 downto 0);
           overread_value : in  STD_LOGIC;
           size : in  STD_LOGIC_VECTOR (1 downto 0);
           connected : in  STD_LOGIC;
           clk : STD_LOGIC);
  end component;

  -- Filtered signals coming from the console
  signal p1_clock_f : std_logic;
  signal p1_latch_f : std_logic;
  signal p2_clock_f : std_logic;
  signal p2_latch_f : std_logic;
  
  -- Toggle signals, useful for monitoring when the FPGA detects a rising edge
  signal p1_clock_toggle : std_logic;
  signal p1_latch_toggle : std_logic;
  signal p1_clock_f_toggle : std_logic;
  signal p1_latch_f_toggle : std_logic;
  signal p2_clock_toggle : std_logic;
  signal p2_latch_toggle : std_logic;
  signal p2_clock_f_toggle : std_logic;
  signal p2_latch_f_toggle : std_logic;
  
  signal data_from_uart : STD_LOGIC_VECTOR (7 downto 0);
  signal uart_data_recieved : STD_LOGIC := '0';
  signal uart_byte_waiting : STD_LOGIC := '0';
  
  signal data_to_uart : STD_LOGIC_VECTOR (7 downto 0) := (others => '0');
  signal uart_buffer_full : STD_LOGIC;
  signal uart_write : STD_LOGIC := '0';
  
  signal serial_receive_mode : std_logic_vector (2 downto 0) := (others => '0');
  signal uart_buffer_ptr : integer range 0 to 16 := 0;
  
  type BUTTON_DATA_buffer is array(0 to 31) of std_logic_vector(31 downto 0);
  
  signal button_queue1 : BUTTON_DATA_BUFFER;
  signal button_queue2 : BUTTON_DATA_BUFFER;
  signal button_queue3 : BUTTON_DATA_BUFFER;
  signal button_queue4 : BUTTON_DATA_BUFFER;
  signal button_queue5 : BUTTON_DATA_BUFFER;
  signal button_queue6 : BUTTON_DATA_BUFFER;
  signal button_queue7 : BUTTON_DATA_BUFFER;
  signal button_queue8 : BUTTON_DATA_BUFFER;
    
  signal buffer_tail : integer range 0 to 31 := 0;
  signal buffer_head : integer range 0 to 31 := 0;
  
  signal prev_latch : std_logic := '0';
  
  signal frame_timer_active : std_logic := '0';
  signal frame_timer : integer range 0 to 160000 := 0;
  
  signal windowed_mode : std_logic := '0';
  
  signal uart_data_temp : std_logic_vector(7 downto 0);
    
  signal controller1_data : std_logic_vector(31 downto 0) := (others => '1');
  signal controller2_data : std_logic_vector(31 downto 0) := (others => '1');
  signal controller3_data : std_logic_vector(31 downto 0) := (others => '1');
  signal controller4_data : std_logic_vector(31 downto 0) := (others => '1');
  signal controller5_data : std_logic_vector(31 downto 0) := (others => '1');
  signal controller6_data : std_logic_vector(31 downto 0) := (others => '1');
  signal controller7_data : std_logic_vector(31 downto 0) := (others => '1');
  signal controller8_data : std_logic_vector(31 downto 0) := (others => '1');
  
  signal controller_size : std_logic_vector(1 downto 0) := "00";
  
  signal controller1_connected : std_logic := '0';
  signal controller2_connected : std_logic := '0';
  signal controller3_connected : std_logic := '0';
  signal controller4_connected : std_logic := '0';
  signal controller5_connected : std_logic := '0';
  signal controller6_connected : std_logic := '0';
  signal controller7_connected : std_logic := '0';
  signal controller8_connected : std_logic := '0';
  
  signal controller1_d0 : std_logic;
  signal controller1_d1 : std_logic;
  signal controller2_d0 : std_logic;
  signal controller2_d1 : std_logic;
  signal controller3_d0 : std_logic;
  signal controller3_d1 : std_logic;
  signal controller4_d0 : std_logic;
  signal controller4_d1 : std_logic;
  signal controller5_d0 : std_logic;
  signal controller5_d1 : std_logic;
  signal controller6_d0 : std_logic;
  signal controller6_d1 : std_logic;
  signal controller7_d0 : std_logic;
  signal controller7_d1 : std_logic;
  signal controller8_d0 : std_logic;
  signal controller8_d1 : std_logic;
  
  signal controller1_d0_oe : std_logic;
  signal controller1_d1_oe : std_logic;
  signal controller2_d0_oe : std_logic;
  signal controller2_d1_oe : std_logic;
  signal controller3_d0_oe : std_logic;
  signal controller3_d1_oe : std_logic;
  signal controller4_d0_oe : std_logic;
  signal controller4_d1_oe : std_logic;
  signal controller5_d0_oe : std_logic;
  signal controller5_d1_oe : std_logic;
  signal controller6_d0_oe : std_logic;
  signal controller6_d1_oe : std_logic;
  signal controller7_d0_oe : std_logic;
  signal controller7_d1_oe : std_logic;
  signal controller8_d0_oe : std_logic;
  signal controller8_d1_oe : std_logic;
begin

  p1_latch_filter: filter port map (signal_in => p1_latch,
                                    clk => CLK,
                                    signal_out => p1_latch_f);
                                 
  p1_clock_filter: filter port map (signal_in => p1_clock,
                                    clk => CLK,
                                    signal_out => p1_clock_f);
                                 
  p2_latch_filter: filter port map (signal_in => p2_latch,
                                    clk => CLK,
                                    signal_out => p2_latch_f);
                                 
  p2_clock_filter: filter port map (signal_in => p2_clock,
                                    clk => CLK,
                                    signal_out => p2_clock_f);
                                    
  p1latch_toggle: toggle port map (signal_in => p1_latch,
                                   signal_out => p1_latch_toggle);
                                 
  p1latch_f_toggle: toggle port map (signal_in => p1_latch_f,
                                     signal_out => p1_latch_f_toggle);
  
  p1clk_toggle: toggle port map (signal_in => p1_clock,
                                 signal_out => p1_clock_toggle);
  
  p1clock_f_toggle: toggle port map (signal_in => p1_clock_f,
                                     signal_out => p1_clock_f_toggle);

  p2latch_toggle: toggle port map (signal_in => p2_latch,
                                   signal_out => p2_latch_toggle);
                                 
  p2latch_f_toggle: toggle port map (signal_in => p2_latch_f,
                                     signal_out => p2_latch_f_toggle);
  
  p2clk_toggle: toggle port map (signal_in => p2_clock,
                                 signal_out => p2_clock_toggle);
  
  p2clock_f_toggle: toggle port map (signal_in => p2_clock_f,
                                     signal_out => p2_clock_f_toggle);
                                     
  uart1: UART port map (rx_data_out => data_from_uart,
                        rx_data_was_recieved => uart_data_recieved,
                        rx_byte_waiting => uart_byte_waiting,
                        clk => CLK,
                        rx_in => RX,
                        tx_data_in => data_to_uart,
                        tx_buffer_full => uart_buffer_full,
                        tx_write => uart_write,
                        tx_out => TX);
                        
  controller1: controller port map (console_clock => p1_clock_f,
                                    console_latch => p1_latch_f,
                                    console_io => '1',
                                    console_d0 => controller1_d0,
                                    console_d1 => controller1_d1,
                                    console_d0_oe => controller1_d0_oe,
                                    console_d1_oe => controller1_d1_oe,
                                    data => controller1_data,
                                    overread_value => '1',
                                    size => controller_size,
                                    connected => controller1_connected,
                                    clk => clk);
                                    
  controller2: controller port map (console_clock => p2_clock_f,
                                    console_latch => p2_latch_f,
                                    console_io => '1',
                                    console_d0 => controller2_d0,
                                    console_d1 => controller2_d1,
                                    console_d0_oe => controller2_d0_oe,
                                    console_d1_oe => controller2_d1_oe,
                                    data => controller2_data,
                                    overread_value => '1',
                                    size => controller_size,
                                    connected => controller2_connected,
                                    clk => clk);
  
  controller3: controller port map (console_clock => p2_clock_f,
                                    console_latch => p2_latch_f,
                                    console_io => '1',
                                    console_d0 => controller3_d0,
                                    console_d1 => controller3_d1,
                                    console_d0_oe => controller3_d0_oe,
                                    console_d1_oe => controller3_d1_oe,
                                    data => controller3_data,
                                    overread_value => '1',
                                    size => controller_size,
                                    connected => controller3_connected,
                                    clk => clk);
  
  controller4: controller port map (console_clock => p2_clock_f,
                                    console_latch => p2_latch_f,
                                    console_io => '1',
                                    console_d0 => controller4_d0,
                                    console_d1 => controller4_d1,
                                    console_d0_oe => controller4_d0_oe,
                                    console_d1_oe => controller4_d1_oe,
                                    data => controller4_data,
                                    overread_value => '1',
                                    size => controller_size,
                                    connected => controller4_connected,
                                    clk => clk);
  
  controller5: controller port map (console_clock => p2_clock_f,
                                    console_latch => p2_latch_f,
                                    console_io => '1',
                                    console_d0 => controller5_d0,
                                    console_d1 => controller5_d1,
                                    console_d0_oe => controller5_d0_oe,
                                    console_d1_oe => controller5_d1_oe,
                                    data => controller5_data,
                                    overread_value => '1',
                                    size => controller_size,
                                    connected => controller5_connected,
                                    clk => clk);  

  controller6: controller port map (console_clock => p2_clock_f,
                                    console_latch => p2_latch_f,
                                    console_io => '1',
                                    console_d0 => controller6_d0,
                                    console_d1 => controller6_d1,
                                    console_d0_oe => controller6_d0_oe,
                                    console_d1_oe => controller6_d1_oe,
                                    data => controller6_data,
                                    overread_value => '1',
                                    size => controller_size,
                                    connected => controller6_connected,
                                    clk => clk); 

  controller7: controller port map (console_clock => p2_clock_f,
                                    console_latch => p2_latch_f,
                                    console_io => '1',
                                    console_d0 => controller7_d0,
                                    console_d1 => controller7_d1,
                                    console_d0_oe => controller7_d0_oe,
                                    console_d1_oe => controller7_d1_oe,
                                    data => controller7_data,
                                    overread_value => '1',
                                    size => controller_size,
                                    connected => controller7_connected,
                                    clk => clk);

  controller8: controller port map (console_clock => p2_clock_f,
                                    console_latch => p2_latch_f,
                                    console_io => '1',
                                    console_d0 => controller8_d0,
                                    console_d1 => controller8_d1,
                                    console_d0_oe => controller8_d0_oe,
                                    console_d1_oe => controller8_d1_oe,
                                    data => controller8_data,
                                    overread_value => '1',
                                    size => controller_size,
                                    connected => controller8_connected,
                                    clk => clk);
                                    
uart_recieve_btye: process(CLK)
	begin
		if (rising_edge(CLK)) then
			if (uart_byte_waiting = '1' and uart_data_recieved = '0') then
        case uart_buffer_ptr is
          when 0 =>
            case data_from_uart is
              when x"66" => -- 'f'
                
                uart_buffer_ptr <= 1;
                serial_receive_mode <= "000";
              
              when x"63" => -- 'c'
                buffer_head <= buffer_tail;
                
                uart_buffer_ptr <= 0;  
              
              when x"77" => -- 'w'
                windowed_mode <= '1';
                
              when x"6C" => -- 'l'
                windowed_mode <= '0';
              
              when x"6E" => -- 'n'
                controller_size <= "00";
                uart_buffer_ptr <= 1;
                serial_receive_mode <= "001";
              
              when x"73" => -- 's'
                controller_size <= "01";
                uart_buffer_ptr <= 1;
                serial_receive_mode <= "010";
              
              when others =>
              
            end case;
            
          when 1 =>
            case serial_receive_mode is
              when "000" =>
                if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
                  button_queue1(buffer_head) <= "111111111111111111111111" & data_from_uart;
                end if;
                
                uart_buffer_ptr <= 2;
              
              when "001" =>
                case data_from_uart is
                  when x"30" => -- '0'
                    controller1_connected <= '0';
                    controller2_connected <= '0';
                    controller3_connected <= '0';
                    controller4_connected <= '0';
                    controller5_connected <= '0';
                    controller6_connected <= '0';
                    controller7_connected <= '0';
                    controller8_connected <= '0';
                  
                  when x"31" => -- '1'
                    controller1_connected <= '1';
                    controller2_connected <= '0';
                    controller3_connected <= '0';
                    controller4_connected <= '0';
                    controller5_connected <= '0';
                    controller6_connected <= '0';
                    controller7_connected <= '0';
                    controller8_connected <= '0';

                  when x"32" => -- '2'
                    controller1_connected <= '1';
                    controller2_connected <= '1';
                    controller3_connected <= '0';
                    controller4_connected <= '0';
                    controller5_connected <= '0';
                    controller6_connected <= '0';
                    controller7_connected <= '0';
                    controller8_connected <= '0';
                  
                  when others =>
                  
                end case;
                
                uart_buffer_ptr <= 0;

              when "010" =>
                case data_from_uart is
                  when x"30" => -- '0'
                    controller1_connected <= '0';
                    controller2_connected <= '0';
                    controller3_connected <= '0';
                    controller4_connected <= '0';
                    controller5_connected <= '0';
                    controller6_connected <= '0';
                    controller7_connected <= '0';
                    controller8_connected <= '0';
                  
                  when x"31" => -- '1'
                    controller1_connected <= '1';
                    controller2_connected <= '0';
                    controller3_connected <= '0';
                    controller4_connected <= '0';
                    controller5_connected <= '0';
                    controller6_connected <= '0';
                    controller7_connected <= '0';
                    controller8_connected <= '0';

                  when x"32" => -- '2'
                    controller1_connected <= '1';
                    controller2_connected <= '1';
                    controller3_connected <= '0';
                    controller4_connected <= '0';
                    controller5_connected <= '0';
                    controller6_connected <= '0';
                    controller7_connected <= '0';
                    controller8_connected <= '0';
                    
                  when x"38" => -- '8'
                    controller1_connected <= '1';
                    controller2_connected <= '1';
                    controller3_connected <= '1';
                    controller4_connected <= '1';
                    controller5_connected <= '1';
                    controller6_connected <= '1';
                    controller7_connected <= '1';
                    controller8_connected <= '1';
                  
                  when others =>
                  
                end case;
                
                uart_buffer_ptr <= 0;
              
              when others =>
                uart_buffer_ptr <= 0;
                
            end case;
            
          when 2 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              if (controller_size = "00") then
                -- add it to the next spot
                button_queue2(buffer_head) <= "111111111111111111111111" & data_from_uart;
                -- move
                if (buffer_head = 31) then
                  buffer_head <= 0;
                else
                  buffer_head <= buffer_head + 1;
                end if;
                uart_buffer_ptr <= 0;
                
              elsif (controller_size = "01") then
                button_queue1(buffer_head) <= "1111111111111111" & data_from_uart & button_queue1(buffer_head)(7 downto 0);
                uart_buffer_ptr <= 3;
              else
                uart_buffer_ptr <= 0;
              end if;
            end if;
            
          when 3 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue2(buffer_head) <= "111111111111111111111111" & data_from_uart;
            end if;  
            uart_buffer_ptr <= 4;
          
          when 4 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue2(buffer_head) <= "1111111111111111" & data_from_uart & button_queue2(buffer_head)(7 downto 0);
            end if;  
            uart_buffer_ptr <= 5;

          when 5 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue3(buffer_head) <= "111111111111111111111111" & data_from_uart;
            end if;  
            uart_buffer_ptr <= 6;
          
          when 6 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue3(buffer_head) <= "1111111111111111" & data_from_uart & button_queue3(buffer_head)(7 downto 0);
            end if;  
            uart_buffer_ptr <= 7;
          
          when 7 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue4(buffer_head) <= "111111111111111111111111" & data_from_uart;
            end if;  
            uart_buffer_ptr <= 8;
          
          when 8 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue4(buffer_head) <= "1111111111111111" & data_from_uart & button_queue4(buffer_head)(7 downto 0);
            end if;  
            uart_buffer_ptr <= 9;

          when 9 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue5(buffer_head) <= "111111111111111111111111" & data_from_uart;
            end if;  
            uart_buffer_ptr <= 10;
          
          when 10 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue5(buffer_head) <= "1111111111111111" & data_from_uart & button_queue5(buffer_head)(7 downto 0);
            end if;  
            uart_buffer_ptr <= 11;
          
          when 11 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue6(buffer_head) <= "111111111111111111111111" & data_from_uart;
            end if;  
            uart_buffer_ptr <= 12;
          
          when 12 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue6(buffer_head) <= "1111111111111111" & data_from_uart & button_queue6(buffer_head)(7 downto 0);
            end if;  
            uart_buffer_ptr <= 13;

          when 13 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue7(buffer_head) <= "111111111111111111111111" & data_from_uart;
            end if;  
            uart_buffer_ptr <= 14;
          
          when 14 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue7(buffer_head) <= "1111111111111111" & data_from_uart & button_queue7(buffer_head)(7 downto 0);
            end if;  
            uart_buffer_ptr <= 15;
          
          when 15 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue8(buffer_head) <= "111111111111111111111111" & data_from_uart;
            end if;  
            uart_buffer_ptr <= 16;
          
          when 16 =>
            if ((buffer_head = 31 and buffer_tail /= 0) or (buffer_head /= 31 and (buffer_head + 1) /= buffer_tail)) then
              button_queue8(buffer_head) <= "1111111111111111" & data_from_uart & button_queue8(buffer_head)(7 downto 0);
              
              -- move
              if (buffer_head = 31) then
                buffer_head <= 0;
              else
                buffer_head <= buffer_head + 1;
              end if;
              uart_buffer_ptr <= 0;              
            end if;  
            uart_buffer_ptr <= 0;
          
          when others =>
        end case;
      	uart_data_recieved <= '1';
			else
				uart_data_recieved <= '0';
			end if;
    end if;
	end process;
  
  process (clk) is
  begin
    if (rising_edge(clk)) then
      uart_write <= '0';
      
      if (windowed_mode = '1' and frame_timer_active = '1') then
        if (frame_timer = 96000) then
          frame_timer <= 0;
          frame_timer_active <= '0';
        
          -- move tail pointer if possible
          if (buffer_tail /= buffer_head) then
            if (buffer_tail = 31) then
              buffer_tail <= 0;
            else
              buffer_tail <= buffer_tail + 1;
            end if;
          end if;
          
          -- Send feedback that a frame was consumed
          if (uart_buffer_full = '0') then
            uart_write <= '1';
            data_to_uart <= x"66";
          end if;
          
        else
          frame_timer <= frame_timer + 1;
        end if;
      end if;

      if (p1_latch_f /= prev_latch) then
        if (p1_latch_f = '1') then
          if (windowed_mode = '1') then
            frame_timer <= 0;
            frame_timer_active <= '1';
          else
            -- move tail pointer if possible
            if (buffer_tail /= buffer_head) then
              if (buffer_tail = 31) then
                buffer_tail <= 0;
              else
                buffer_tail <= buffer_tail + 1;
              end if;
            end if;
            
            -- Send feedback that a frame was consumed
            if (uart_buffer_full = '0') then
              uart_write <= '1';
              data_to_uart <= x"66";
            end if;
          end if;
        end if;
        prev_latch <= p1_latch_f;
      end if;
    end if;
  end process;

  controller1_data <= button_queue1(buffer_tail) when buffer_head /= buffer_tail else
                      button_queue1(31) when buffer_tail = 0 else
                      button_queue1(buffer_tail-1);

  controller2_data <= button_queue2(buffer_tail) when buffer_head /= buffer_tail else
                      button_queue2(31) when buffer_tail = 0 else
                      button_queue2(buffer_tail-1);
  
  controller3_data <= button_queue3(buffer_tail) when buffer_head /= buffer_tail else
                      button_queue3(31) when buffer_tail = 0 else
                      button_queue3(buffer_tail-1);

  controller4_data <= button_queue4(buffer_tail) when buffer_head /= buffer_tail else
                      button_queue4(31) when buffer_tail = 0 else
                      button_queue4(buffer_tail-1);
                      
  controller5_data <= button_queue5(buffer_tail) when buffer_head /= buffer_tail else
                      button_queue5(31) when buffer_tail = 0 else
                      button_queue5(buffer_tail-1);

  controller6_data <= button_queue6(buffer_tail) when buffer_head /= buffer_tail else
                      button_queue6(31) when buffer_tail = 0 else
                      button_queue6(buffer_tail-1);
                      
  controller7_data <= button_queue7(buffer_tail) when buffer_head /= buffer_tail else
                      button_queue7(31) when buffer_tail = 0 else
                      button_queue7(buffer_tail-1);

  controller8_data <= button_queue8(buffer_tail) when buffer_head /= buffer_tail else
                      button_queue8(31) when buffer_tail = 0 else
                      button_queue8(buffer_tail-1);

  p1_d0 <= controller1_d0;
  p1_d1 <= controller1_d1;
  p2_d0 <= controller2_d0;
  p2_d1 <= controller2_d1;
  
  p1_d0_oe <= controller1_d0_oe;
  p1_d1_oe <= controller1_d1_oe;
  p2_d0_oe <= controller2_d0_oe;
  p2_d1_oe <= controller2_d1_oe;
  

  l <= std_logic_vector(to_unsigned(buffer_tail, 4));
    
  debug(0) <= p1_latch_toggle;
  debug(1) <= p2_latch_f;
  debug(2) <= p1_clock_toggle;
  debug(3) <= p2_clock_f;

end Behavioral;

